module layer2_rom (
    output signed [7:0] w0_0,
    output signed [7:0] w0_1,
    output signed [7:0] w0_2,
    output signed [7:0] w0_3,
    output signed [7:0] w0_4,
    output signed [7:0] w0_5,
    output signed [7:0] w0_6,
    output signed [7:0] w0_7,
    output signed [7:0] w1_0,
    output signed [7:0] w1_1,
    output signed [7:0] w1_2,
    output signed [7:0] w1_3,
    output signed [7:0] w1_4,
    output signed [7:0] w1_5,
    output signed [7:0] w1_6,
    output signed [7:0] w1_7,
    output signed [7:0] w2_0,
    output signed [7:0] w2_1,
    output signed [7:0] w2_2,
    output signed [7:0] w2_3,
    output signed [7:0] w2_4,
    output signed [7:0] w2_5,
    output signed [7:0] w2_6,
    output signed [7:0] w2_7,
    output signed [7:0] w3_0,
    output signed [7:0] w3_1,
    output signed [7:0] w3_2,
    output signed [7:0] w3_3,
    output signed [7:0] w3_4,
    output signed [7:0] w3_5,
    output signed [7:0] w3_6,
    output signed [7:0] w3_7,
    output signed [7:0] w4_0,
    output signed [7:0] w4_1,
    output signed [7:0] w4_2,
    output signed [7:0] w4_3,
    output signed [7:0] w4_4,
    output signed [7:0] w4_5,
    output signed [7:0] w4_6,
    output signed [7:0] w4_7,
    output signed [7:0] w5_0,
    output signed [7:0] w5_1,
    output signed [7:0] w5_2,
    output signed [7:0] w5_3,
    output signed [7:0] w5_4,
    output signed [7:0] w5_5,
    output signed [7:0] w5_6,
    output signed [7:0] w5_7,
    output signed [7:0] w6_0,
    output signed [7:0] w6_1,
    output signed [7:0] w6_2,
    output signed [7:0] w6_3,
    output signed [7:0] w6_4,
    output signed [7:0] w6_5,
    output signed [7:0] w6_6,
    output signed [7:0] w6_7,
    output signed [7:0] w7_0,
    output signed [7:0] w7_1,
    output signed [7:0] w7_2,
    output signed [7:0] w7_3,
    output signed [7:0] w7_4,
    output signed [7:0] w7_5,
    output signed [7:0] w7_6,
    output signed [7:0] w7_7,
    output signed [7:0] b0,
    output signed [7:0] b1,
    output signed [7:0] b2,
    output signed [7:0] b3,
    output signed [7:0] b4,
    output signed [7:0] b5,
    output signed [7:0] b6,
    output signed [7:0] b7
);

    // Auto-generated from trained model

    assign w0_0 = -76;
    assign w0_1 = 4;
    assign w0_2 = -28;
    assign w0_3 = 14;
    assign w0_4 = -71;
    assign w0_5 = -40;
    assign w0_6 = -38;
    assign w0_7 = -35;
    assign w1_0 = -38;
    assign w1_1 = 3;
    assign w1_2 = -25;
    assign w1_3 = 11;
    assign w1_4 = -32;
    assign w1_5 = -26;
    assign w1_6 = -22;
    assign w1_7 = -27;
    assign w2_0 = -47;
    assign w2_1 = 4;
    assign w2_2 = -23;
    assign w2_3 = 9;
    assign w2_4 = -45;
    assign w2_5 = -25;
    assign w2_6 = -23;
    assign w2_7 = -21;
    assign w3_0 = 8;
    assign w3_1 = 32;
    assign w3_2 = 77;
    assign w3_3 = -1;
    assign w3_4 = 9;
    assign w3_5 = 3;
    assign w3_6 = 83;
    assign w3_7 = 72;
    assign w4_0 = -2;
    assign w4_1 = -30;
    assign w4_2 = -72;
    assign w4_3 = -53;
    assign w4_4 = 127;
    assign w4_5 = 2;
    assign w4_6 = -35;
    assign w4_7 = -24;
    assign w5_0 = -3;
    assign w5_1 = 25;
    assign w5_2 = 29;
    assign w5_3 = 84;
    assign w5_4 = -1;
    assign w5_5 = -1;
    assign w5_6 = 33;
    assign w5_7 = 9;
    assign w6_0 = 32;
    assign w6_1 = -32;
    assign w6_2 = 2;
    assign w6_3 = -10;
    assign w6_4 = 12;
    assign w6_5 = 29;
    assign w6_6 = 6;
    assign w6_7 = -49;
    assign w7_0 = -4;
    assign w7_1 = -8;
    assign w7_2 = 42;
    assign w7_3 = 1;
    assign w7_4 = 0;
    assign w7_5 = -5;
    assign w7_6 = 43;
    assign w7_7 = 82;
    assign b0 = 29;
    assign b1 = -72;
    assign b2 = 22;
    assign b3 = 119;
    assign b4 = 5;
    assign b5 = -127;
    assign b6 = 39;
    assign b7 = 41;
endmodule
