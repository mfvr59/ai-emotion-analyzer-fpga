module layer1_rom (
    output signed [7:0] w0_0,
    output signed [7:0] w0_1,
    output signed [7:0] w0_2,
    output signed [7:0] w0_3,
    output signed [7:0] w0_4,
    output signed [7:0] w0_5,
    output signed [7:0] w0_6,
    output signed [7:0] w0_7,
    output signed [7:0] w0_8,
    output signed [7:0] w0_9,
    output signed [7:0] w0_10,
    output signed [7:0] w0_11,
    output signed [7:0] w0_12,
    output signed [7:0] w0_13,
    output signed [7:0] w0_14,
    output signed [7:0] w0_15,
    output signed [7:0] w1_0,
    output signed [7:0] w1_1,
    output signed [7:0] w1_2,
    output signed [7:0] w1_3,
    output signed [7:0] w1_4,
    output signed [7:0] w1_5,
    output signed [7:0] w1_6,
    output signed [7:0] w1_7,
    output signed [7:0] w1_8,
    output signed [7:0] w1_9,
    output signed [7:0] w1_10,
    output signed [7:0] w1_11,
    output signed [7:0] w1_12,
    output signed [7:0] w1_13,
    output signed [7:0] w1_14,
    output signed [7:0] w1_15,
    output signed [7:0] w2_0,
    output signed [7:0] w2_1,
    output signed [7:0] w2_2,
    output signed [7:0] w2_3,
    output signed [7:0] w2_4,
    output signed [7:0] w2_5,
    output signed [7:0] w2_6,
    output signed [7:0] w2_7,
    output signed [7:0] w2_8,
    output signed [7:0] w2_9,
    output signed [7:0] w2_10,
    output signed [7:0] w2_11,
    output signed [7:0] w2_12,
    output signed [7:0] w2_13,
    output signed [7:0] w2_14,
    output signed [7:0] w2_15,
    output signed [7:0] w3_0,
    output signed [7:0] w3_1,
    output signed [7:0] w3_2,
    output signed [7:0] w3_3,
    output signed [7:0] w3_4,
    output signed [7:0] w3_5,
    output signed [7:0] w3_6,
    output signed [7:0] w3_7,
    output signed [7:0] w3_8,
    output signed [7:0] w3_9,
    output signed [7:0] w3_10,
    output signed [7:0] w3_11,
    output signed [7:0] w3_12,
    output signed [7:0] w3_13,
    output signed [7:0] w3_14,
    output signed [7:0] w3_15,
    output signed [7:0] w4_0,
    output signed [7:0] w4_1,
    output signed [7:0] w4_2,
    output signed [7:0] w4_3,
    output signed [7:0] w4_4,
    output signed [7:0] w4_5,
    output signed [7:0] w4_6,
    output signed [7:0] w4_7,
    output signed [7:0] w4_8,
    output signed [7:0] w4_9,
    output signed [7:0] w4_10,
    output signed [7:0] w4_11,
    output signed [7:0] w4_12,
    output signed [7:0] w4_13,
    output signed [7:0] w4_14,
    output signed [7:0] w4_15,
    output signed [7:0] w5_0,
    output signed [7:0] w5_1,
    output signed [7:0] w5_2,
    output signed [7:0] w5_3,
    output signed [7:0] w5_4,
    output signed [7:0] w5_5,
    output signed [7:0] w5_6,
    output signed [7:0] w5_7,
    output signed [7:0] w5_8,
    output signed [7:0] w5_9,
    output signed [7:0] w5_10,
    output signed [7:0] w5_11,
    output signed [7:0] w5_12,
    output signed [7:0] w5_13,
    output signed [7:0] w5_14,
    output signed [7:0] w5_15,
    output signed [7:0] w6_0,
    output signed [7:0] w6_1,
    output signed [7:0] w6_2,
    output signed [7:0] w6_3,
    output signed [7:0] w6_4,
    output signed [7:0] w6_5,
    output signed [7:0] w6_6,
    output signed [7:0] w6_7,
    output signed [7:0] w6_8,
    output signed [7:0] w6_9,
    output signed [7:0] w6_10,
    output signed [7:0] w6_11,
    output signed [7:0] w6_12,
    output signed [7:0] w6_13,
    output signed [7:0] w6_14,
    output signed [7:0] w6_15,
    output signed [7:0] w7_0,
    output signed [7:0] w7_1,
    output signed [7:0] w7_2,
    output signed [7:0] w7_3,
    output signed [7:0] w7_4,
    output signed [7:0] w7_5,
    output signed [7:0] w7_6,
    output signed [7:0] w7_7,
    output signed [7:0] w7_8,
    output signed [7:0] w7_9,
    output signed [7:0] w7_10,
    output signed [7:0] w7_11,
    output signed [7:0] w7_12,
    output signed [7:0] w7_13,
    output signed [7:0] w7_14,
    output signed [7:0] w7_15,
    output signed [7:0] b0,
    output signed [7:0] b1,
    output signed [7:0] b2,
    output signed [7:0] b3,
    output signed [7:0] b4,
    output signed [7:0] b5,
    output signed [7:0] b6,
    output signed [7:0] b7
);

    // Auto-generated from trained model
    assign w0_0 = -14;
    assign w0_1 = -8;
    assign w0_2 = -25;
    assign w0_3 = -11;
    assign w0_4 = 2;
    assign w0_5 = 15;
    assign w0_6 = 31;
    assign w0_7 = 35;
    assign w0_8 = 36;
    assign w0_9 = -7;
    assign w0_10 = -18;
    assign w0_11 = 8;
    assign w0_12 = -127;
    assign w0_13 = -12;
    assign w0_14 = -29;
    assign w0_15 = 60;
    assign w1_0 = 35;
    assign w1_1 = 35;
    assign w1_2 = -26;
    assign w1_3 = 14;
    assign w1_4 = 19;
    assign w1_5 = -48;
    assign w1_6 = -47;
    assign w1_7 = -79;
    assign w1_8 = -79;
    assign w1_9 = -24;
    assign w1_10 = 9;
    assign w1_11 = -9;
    assign w1_12 = -26;
    assign w1_13 = -9;
    assign w1_14 = 52;
    assign w1_15 = -74;
    assign w2_0 = -4;
    assign w2_1 = 5;
    assign w2_2 = 9;
    assign w2_3 = 13;
    assign w2_4 = 16;
    assign w2_5 = 29;
    assign w2_6 = 59;
    assign w2_7 = 60;
    assign w2_8 = 57;
    assign w2_9 = -13;
    assign w2_10 = -11;
    assign w2_11 = 11;
    assign w2_12 = -5;
    assign w2_13 = -17;
    assign w2_14 = -38;
    assign w2_15 = 80;
    assign w3_0 = 9;
    assign w3_1 = 43;
    assign w3_2 = -7;
    assign w3_3 = 11;
    assign w3_4 = 32;
    assign w3_5 = -33;
    assign w3_6 = -4;
    assign w3_7 = -59;
    assign w3_8 = -55;
    assign w3_9 = 50;
    assign w3_10 = 41;
    assign w3_11 = -34;
    assign w3_12 = -11;
    assign w3_13 = -41;
    assign w3_14 = 12;
    assign w3_15 = -28;
    assign w4_0 = -4;
    assign w4_1 = -35;
    assign w4_2 = -78;
    assign w4_3 = -17;
    assign w4_4 = -10;
    assign w4_5 = 46;
    assign w4_6 = 54;
    assign w4_7 = 69;
    assign w4_8 = 65;
    assign w4_9 = 15;
    assign w4_10 = -33;
    assign w4_11 = 21;
    assign w4_12 = -28;
    assign w4_13 = 8;
    assign w4_14 = -49;
    assign w4_15 = 28;
    assign w5_0 = -63;
    assign w5_1 = 4;
    assign w5_2 = -38;
    assign w5_3 = -51;
    assign w5_4 = -40;
    assign w5_5 = -70;
    assign w5_6 = 31;
    assign w5_7 = -53;
    assign w5_8 = -29;
    assign w5_9 = -28;
    assign w5_10 = 18;
    assign w5_11 = 27;
    assign w5_12 = 12;
    assign w5_13 = -52;
    assign w5_14 = -49;
    assign w5_15 = -46;
    assign w6_0 = -54;
    assign w6_1 = -40;
    assign w6_2 = 7;
    assign w6_3 = -28;
    assign w6_4 = -12;
    assign w6_5 = 42;
    assign w6_6 = 36;
    assign w6_7 = 86;
    assign w6_8 = 83;
    assign w6_9 = 54;
    assign w6_10 = 37;
    assign w6_11 = 33;
    assign w6_12 = 37;
    assign w6_13 = 34;
    assign w6_14 = 14;
    assign w6_15 = 59;
    assign w7_0 = 26;
    assign w7_1 = -6;
    assign w7_2 = 3;
    assign w7_3 = -2;
    assign w7_4 = -26;
    assign w7_5 = -58;
    assign w7_6 = -71;
    assign w7_7 = -80;
    assign w7_8 = -76;
    assign w7_9 = -21;
    assign w7_10 = -1;
    assign w7_11 = -9;
    assign w7_12 = 22;
    assign w7_13 = 16;
    assign w7_14 = 33;
    assign w7_15 = -82;
    assign b0 = -50;
    assign b1 = 73;
    assign b2 = 97;
    assign b3 = -100;
    assign b4 = 63;
    assign b5 = -44;
    assign b6 = 7;
    assign b7 = 127;
endmodule
