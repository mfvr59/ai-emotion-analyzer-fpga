module layer3_rom (
    output signed [7:0] w0_0,
    output signed [7:0] w0_1,
    output signed [7:0] w0_2,
    output signed [7:0] w0_3,
    output signed [7:0] w0_4,
    output signed [7:0] w0_5,
    output signed [7:0] w0_6,
    output signed [7:0] w0_7,
    output signed [7:0] w1_0,
    output signed [7:0] w1_1,
    output signed [7:0] w1_2,
    output signed [7:0] w1_3,
    output signed [7:0] w1_4,
    output signed [7:0] w1_5,
    output signed [7:0] w1_6,
    output signed [7:0] w1_7,
    output signed [7:0] w2_0,
    output signed [7:0] w2_1,
    output signed [7:0] w2_2,
    output signed [7:0] w2_3,
    output signed [7:0] w2_4,
    output signed [7:0] w2_5,
    output signed [7:0] w2_6,
    output signed [7:0] w2_7,
    output signed [7:0] w3_0,
    output signed [7:0] w3_1,
    output signed [7:0] w3_2,
    output signed [7:0] w3_3,
    output signed [7:0] w3_4,
    output signed [7:0] w3_5,
    output signed [7:0] w3_6,
    output signed [7:0] w3_7,
    output signed [7:0] w4_0,
    output signed [7:0] w4_1,
    output signed [7:0] w4_2,
    output signed [7:0] w4_3,
    output signed [7:0] w4_4,
    output signed [7:0] w4_5,
    output signed [7:0] w4_6,
    output signed [7:0] w4_7,
    output signed [7:0] w5_0,
    output signed [7:0] w5_1,
    output signed [7:0] w5_2,
    output signed [7:0] w5_3,
    output signed [7:0] w5_4,
    output signed [7:0] w5_5,
    output signed [7:0] w5_6,
    output signed [7:0] w5_7,
    output signed [7:0] w6_0,
    output signed [7:0] w6_1,
    output signed [7:0] w6_2,
    output signed [7:0] w6_3,
    output signed [7:0] w6_4,
    output signed [7:0] w6_5,
    output signed [7:0] w6_6,
    output signed [7:0] w6_7,
    output signed [7:0] w7_0,
    output signed [7:0] w7_1,
    output signed [7:0] w7_2,
    output signed [7:0] w7_3,
    output signed [7:0] w7_4,
    output signed [7:0] w7_5,
    output signed [7:0] w7_6,
    output signed [7:0] w7_7,
    output signed [7:0] b0,
    output signed [7:0] b1,
    output signed [7:0] b2,
    output signed [7:0] b3,
    output signed [7:0] b4,
    output signed [7:0] b5,
    output signed [7:0] b6,
    output signed [7:0] b7
);

    // Auto-generated from trained model
    assign w0_0 = 63;
    assign w0_1 = 46;
    assign w0_2 = 72;
    assign w0_3 = -22;
    assign w0_4 = -127;
    assign w0_5 = 27;
    assign w0_6 = -87;
    assign w0_7 = 2;
    assign w1_0 = -45;
    assign w1_1 = -46;
    assign w1_2 = -10;
    assign w1_3 = -67;
    assign w1_4 = 19;
    assign w1_5 = -127;
    assign w1_6 = 19;
    assign w1_7 = -48;
    assign w2_0 = -29;
    assign w2_1 = -16;
    assign w2_2 = 3;
    assign w2_3 = 61;
    assign w2_4 = -18;
    assign w2_5 = 26;
    assign w2_6 = 10;
    assign w2_7 = 46;
    assign w3_0 = 0;
    assign w3_1 = 0;
    assign w3_2 = 0;
    assign w3_3 = 0;
    assign w3_4 = 0;
    assign w3_5 = 0;
    assign w3_6 = 0;
    assign w3_7 = 0;
    assign w4_0 = 0;
    assign w4_1 = 0;
    assign w4_2 = 0;
    assign w4_3 = 0;
    assign w4_4 = 0;
    assign w4_5 = 0;
    assign w4_6 = 0;
    assign w4_7 = 0;
    assign w5_0 = 0;
    assign w5_1 = 0;
    assign w5_2 = 0;
    assign w5_3 = 0;
    assign w5_4 = 0;
    assign w5_5 = 0;
    assign w5_6 = 0;
    assign w5_7 = 0;
    assign w6_0 = 0;
    assign w6_1 = 0;
    assign w6_2 = 0;
    assign w6_3 = 0;
    assign w6_4 = 0;
    assign w6_5 = 0;
    assign w6_6 = 0;
    assign w6_7 = 0;
    assign w7_0 = 0;
    assign w7_1 = 0;
    assign w7_2 = 0;
    assign w7_3 = 0;
    assign w7_4 = 0;
    assign w7_5 = 0;
    assign w7_6 = 0;
    assign w7_7 = 0;
    assign b0 = -75;
    assign b1 = 127;
    assign b2 = -20; 
    assign b3 = 0; 
    assign b4 = 0;
    assign b5 = 0; 
    assign b6 = 0;
    assign b7 = 0;
endmodule
